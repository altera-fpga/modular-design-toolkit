/* ##################################################################################
�* Copyright (C) 2025 Intel Corporation
 *
�* This software and the related documents are Intel copyrighted materials, and
 * your use of them is governed by the express license under which they were
 * provided to you ("License"). Unless the License provides otherwise, you may
 * not use, modify, copy, publish, distribute, disclose or transmit this software
 * or the related documents without Intel's prior written permission.
 *
�* This software and the related documents are provided as is, with no express
�* or implied warranties, other than those that are expressly stated in the License.
 * ##################################################################################

 * ##################################################################################
 *
 * Module: intel_vvp_reset_extend
 *
 * Description: extends reset duration
 *
 * ##################################################################################
*/

`default_nettype none

module intel_issp_reset_shim (
  issp_in,
  reset_out
);

  input    wire    issp_in;
  output   wire    reset_out;

  assign reset_out  = issp_in;

endmodule

`default_nettype wire
